module tb;
    
    initial begin
        $system("mv design.v adder.v")
    end

endmodule : tb