always @(posedge clk or negedge reset) begin
    if(~reset)
end

always @(posedge clk) begin
    if(~reset)
end