package sfr_pkg;
    `include "sfr_item.sv"
    `include "reg2sfr_adapter.sv"
    `include "sfr_master_monitor.sv"
    `include "sfr_master_driver.sv"
    `include "sfr_master_sequencer.sv"
    `include "sfr_master_agent.sv"
endpackage : sfr_pkg